<?xml version="1.0" encoding="UTF-8"?>
<Batch version="2.0"><TaskList><Task type="CropTask" enabled="True"><Left units="0" base_point="0">0</Left><Right units="0" base_point="0">1545</Right><Top units="0" base_point="0">0</Top><Bottom units="0" base_point="2">0</Bottom><Color>#FFFFFF</Color><Alpha>255</Alpha><BlurredImage>False</BlurredImage></Task><Task type="ResizeTask" enabled="True"><Width units="0">500</Width><Height units="0">-1</Height><DPI>-1</DPI><Filter>9</Filter><UseProportions>True</UseProportions><ResizeType>0</ResizeType></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>_Back]]></FileName><PreserveStruct>False</PreserveStruct><CommonFolder><![CDATA[C:\Users\krobison\Downloads\]]></CommonFolder><FileType>JPG</FileType><FilePath><![CDATA[<Source Folder>]]></FilePath><FileExists>0</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed><DDSMIPLevels>8</DDSMIPLevels><DDSMipMapFilter>4</DDSMipMapFilter><DDSFormat>71</DDSFormat></Task></TaskList></Batch>
